module clock_gen (
    output logic clock
);
    
endmodule