module commutator (
    ports
);
    
endmodule