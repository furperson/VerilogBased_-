module control_unit (
    ports
);
    
endmodule