module ALU (
    input logic [15:0] argA_i,
    input logic [15:0] argB_i,
    input logic isInvertA_i,
    input logic isInvertB_i,
    input logic isInc_i,
    input logic isAnd_i
    output logic result_o,
);
    
endmodule